module top(
    input [6:0]sw,
    output [1:0]led
);

endmodule
